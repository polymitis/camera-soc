// Project : camera_fpga_app
// Author  : Petros Fountas
// Details : Top module for Terasic DE1-SOC rev.D board.
`include "TRDB_D5M.sv"

module CameraFpga (
    input logic         piul1FpgaClock,
    input logic         piul1FpgaResetn,
    tITRDB_D5M.driver   pIImageSensor
    );



endmodule
